magic
tech scmos
timestamp 1715202207
<< polysilicon >>
rect -15 39 -13 41
rect -7 39 -5 41
rect -15 11 -13 26
rect -7 11 -5 26
rect -15 -1 -13 1
rect -7 -1 -5 1
<< ndiffusion >>
rect -16 1 -15 11
rect -13 1 -7 11
rect -5 1 -4 11
<< pdiffusion >>
rect -16 26 -15 39
rect -13 26 -12 39
rect -8 26 -7 39
rect -5 26 -4 39
<< metal1 >>
rect -20 47 0 48
rect -20 43 -19 47
rect -15 43 -5 47
rect -1 43 0 47
rect -20 42 0 43
rect -20 39 -16 42
rect -4 39 0 42
rect -12 16 -8 26
rect -1 19 0 23
rect -12 12 0 16
rect -4 11 0 12
rect -20 -2 -16 1
rect -20 -3 0 -2
rect -20 -7 -19 -3
rect -15 -7 -5 -3
rect -1 -7 0 -3
rect -20 -8 0 -7
<< ntransistor >>
rect -15 1 -13 11
rect -7 1 -5 11
<< ptransistor >>
rect -15 26 -13 39
rect -7 26 -5 39
<< polycontact >>
rect -19 19 -15 23
rect -5 19 -1 23
<< ndcontact >>
rect -20 1 -16 11
rect -4 1 0 11
<< pdcontact >>
rect -20 26 -16 39
rect -12 26 -8 39
rect -4 26 0 39
<< psubstratepcontact >>
rect -19 -7 -15 -3
rect -5 -7 -1 -3
<< nsubstratencontact >>
rect -19 43 -15 47
rect -5 43 -1 47
<< labels >>
rlabel polycontact -18 21 -18 21 3 IN1
rlabel metal1 -10 47 -10 47 5 VDD
rlabel metal1 -10 -5 -10 -5 1 GND
rlabel metal1 -2 14 -2 14 7 OUT
rlabel polycontact -1 21 -1 21 7 IN2
<< end >>
